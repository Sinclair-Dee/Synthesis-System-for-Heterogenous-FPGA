// megafunction wizard: %ALTMULT_ACCUM (MAC)%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altmult_add 

// ============================================================
// File Name: mult.v
// Megafunction Name(s):
// 			altmult_add
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 13.0.1 Build 232 06/12/2013 SP 1 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2013 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module mult (
	accum_sload,
	aclr3,
	clock0,
	dataa_0,
	dataa_1,
	datab_0,
	datab_1,
	ena0,
	result);

	input	  accum_sload;
	input	  aclr3;
	input	  clock0;
	input	[15:0]  dataa_0;
	input	[15:0]  dataa_1;
	input	[15:0]  datab_0;
	input	[15:0]  datab_1;
	input	  ena0;
	output	[43:0]  result;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri0	  accum_sload;
	tri0	  aclr3;
	tri1	  clock0;
	tri0	[15:0]  dataa_0;
	tri0	[15:0]  dataa_1;
	tri0	[15:0]  datab_0;
	tri0	[15:0]  datab_1;
	tri1	  ena0;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire [43:0] sub_wire0;
	wire [15:0] sub_wire6 = dataa_1[15:0];
	wire [15:0] sub_wire3 = datab_1[15:0];
	wire [43:0] result = sub_wire0[43:0];
	wire [15:0] sub_wire1 = datab_0[15:0];
	wire [31:0] sub_wire2 = {sub_wire3, sub_wire1};
	wire [15:0] sub_wire4 = dataa_0[15:0];
	wire [31:0] sub_wire5 = {sub_wire6, sub_wire4};

	altmult_add	altmult_add_component (
				.clock0 (clock0),
				.datab (sub_wire2),
				.ena0 (ena0),
				.accum_sload (accum_sload),
				.aclr3 (aclr3),
				.dataa (sub_wire5),
				.result (sub_wire0),
				.aclr0 (1'b0),
				.aclr1 (1'b0),
				.aclr2 (1'b0),
				.addnsub1 (1'b1),
				.addnsub1_round (1'b0),
				.addnsub3 (1'b1),
				.addnsub3_round (1'b0),
				.chainin (1'b0),
				.chainout_round (1'b0),
				.chainout_sat_overflow (),
				.chainout_saturate (1'b0),
				.clock1 (1'b1),
				.clock2 (1'b1),
				.clock3 (1'b1),
				.coefsel0 ({3{1'b0}}),
				.coefsel1 ({3{1'b0}}),
				.coefsel2 ({3{1'b0}}),
				.coefsel3 ({3{1'b0}}),
				.datac ({44{1'b0}}),
				.ena1 (1'b1),
				.ena2 (1'b1),
				.ena3 (1'b1),
				.mult01_round (1'b0),
				.mult01_saturation (1'b0),
				.mult0_is_saturated (),
				.mult1_is_saturated (),
				.mult23_round (1'b0),
				.mult23_saturation (1'b0),
				.mult2_is_saturated (),
				.mult3_is_saturated (),
				.output_round (1'b0),
				.output_saturate (1'b0),
				.overflow (),
				.rotate (1'b0),
				.scanina ({16{1'b0}}),
				.scaninb ({16{1'b0}}),
				.scanouta (),
				.scanoutb (),
				.shift_right (1'b0),
				.signa (1'b0),
				.signb (1'b0),
				.sourcea ({2{1'b0}}),
				.sourceb ({2{1'b0}}),
				.zero_chainout (1'b0),
				.zero_loopback (1'b0));
	defparam
		altmult_add_component.accumulator = "YES",
		altmult_add_component.accum_direction = "ADD",
		altmult_add_component.accum_sload_aclr = "ACLR3",
		altmult_add_component.accum_sload_pipeline_aclr = "ACLR3",
		altmult_add_component.accum_sload_pipeline_register = "CLOCK0",
		altmult_add_component.accum_sload_register = "CLOCK0",
		altmult_add_component.addnsub_multiplier_aclr1 = "ACLR3",
		altmult_add_component.addnsub_multiplier_pipeline_aclr1 = "ACLR3",
		altmult_add_component.addnsub_multiplier_pipeline_register1 = "CLOCK0",
		altmult_add_component.addnsub_multiplier_register1 = "CLOCK0",
		altmult_add_component.chainout_adder = "NO",
		altmult_add_component.chainout_register = "UNREGISTERED",
		altmult_add_component.dedicated_multiplier_circuitry = "AUTO",
		altmult_add_component.input_aclr_a0 = "ACLR3",
		altmult_add_component.input_aclr_a1 = "ACLR3",
		altmult_add_component.input_aclr_b0 = "ACLR3",
		altmult_add_component.input_aclr_b1 = "ACLR3",
		altmult_add_component.input_register_a0 = "CLOCK0",
		altmult_add_component.input_register_a1 = "CLOCK0",
		altmult_add_component.input_register_b0 = "CLOCK0",
		altmult_add_component.input_register_b1 = "CLOCK0",
		altmult_add_component.input_source_a0 = "DATAA",
		altmult_add_component.input_source_a1 = "DATAA",
		altmult_add_component.input_source_b0 = "DATAB",
		altmult_add_component.input_source_b1 = "DATAB",
		altmult_add_component.intended_device_family = "Stratix III",
		altmult_add_component.lpm_type = "altmult_add",
		altmult_add_component.multiplier1_direction = "ADD",
		altmult_add_component.multiplier_aclr0 = "ACLR3",
		altmult_add_component.multiplier_aclr1 = "ACLR3",
		altmult_add_component.multiplier_register0 = "CLOCK0",
		altmult_add_component.multiplier_register1 = "CLOCK0",
		altmult_add_component.number_of_multipliers = 2,
		altmult_add_component.output_aclr = "ACLR3",
		altmult_add_component.output_register = "CLOCK0",
		altmult_add_component.port_addnsub1 = "PORT_UNUSED",
		altmult_add_component.port_signa = "PORT_UNUSED",
		altmult_add_component.port_signb = "PORT_UNUSED",
		altmult_add_component.representation_a = "SIGNED",
		altmult_add_component.representation_b = "SIGNED",
		altmult_add_component.signed_aclr_a = "ACLR3",
		altmult_add_component.signed_aclr_b = "ACLR3",
		altmult_add_component.signed_pipeline_aclr_a = "ACLR3",
		altmult_add_component.signed_pipeline_aclr_b = "ACLR3",
		altmult_add_component.signed_pipeline_register_a = "CLOCK0",
		altmult_add_component.signed_pipeline_register_b = "CLOCK0",
		altmult_add_component.signed_register_a = "CLOCK0",
		altmult_add_component.signed_register_b = "CLOCK0",
		altmult_add_component.width_a = 16,
		altmult_add_component.width_b = 16,
		altmult_add_component.width_chainin = 1,
		altmult_add_component.width_result = 44,
		altmult_add_component.zero_chainout_output_register = "UNREGISTERED",
		altmult_add_component.zero_loopback_aclr = "ACLR3",
		altmult_add_component.zero_loopback_output_aclr = "ACLR3",
		altmult_add_component.zero_loopback_output_register = "CLOCK0",
		altmult_add_component.zero_loopback_pipeline_aclr = "ACLR3",
		altmult_add_component.zero_loopback_pipeline_register = "CLOCK0",
		altmult_add_component.zero_loopback_register = "CLOCK0";


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ACCUM_DIRECTION STRING "Add"
// Retrieval info: PRIVATE: ACCUM_SLOAD NUMERIC "1"
// Retrieval info: PRIVATE: ACCUM_SLOAD_ACLR NUMERIC "3"
// Retrieval info: PRIVATE: ACCUM_SLOAD_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ACCUM_SLOAD_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ACCUM_SLOAD_PIPELINE_ACLR NUMERIC "3"
// Retrieval info: PRIVATE: ACCUM_SLOAD_PIPELINE_REG NUMERIC "1"
// Retrieval info: PRIVATE: ACCUM_SLOAD_PIPELINE_REG_INDEX NUMERIC "0"
// Retrieval info: PRIVATE: ACCUM_SLOAD_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ACCUM_SLOAD_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ACCUM_SLOAD_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: ACCUM_SLOAD_REG NUMERIC "1"
// Retrieval info: PRIVATE: ACCUM_SLOAD_REG_INDEX NUMERIC "0"
// Retrieval info: PRIVATE: ACCUM_SLOAD_UPPER_DATA NUMERIC "0"
// Retrieval info: PRIVATE: ACCUM_SLOAD_UPPER_DATA_ACLR NUMERIC "3"
// Retrieval info: PRIVATE: ACCUM_SLOAD_UPPER_DATA_PIPELINE_ACLR NUMERIC "3"
// Retrieval info: PRIVATE: ACCUM_SLOAD_UPPER_DATA_PIPELINE_REG NUMERIC "0"
// Retrieval info: PRIVATE: ACCUM_SLOAD_UPPER_DATA_REG NUMERIC "0"
// Retrieval info: PRIVATE: ADDNSUB1_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ADDNSUB1_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ADDNSUB1_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ADDNSUB1_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ADDNSUB1_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: ADDNSUB1_REG STRING "1"
// Retrieval info: PRIVATE: ADDNSUB3_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ADDNSUB3_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ADDNSUB3_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ADDNSUB3_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ADDNSUB3_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: ADDNSUB3_REG STRING "1"
// Retrieval info: PRIVATE: ADD_ENABLE NUMERIC "1"
// Retrieval info: PRIVATE: ALL_REG_ACLR NUMERIC "1"
// Retrieval info: PRIVATE: A_ACLR_SRC_MULT0 NUMERIC "3"
// Retrieval info: PRIVATE: A_CLK_SRC_MULT0 NUMERIC "0"
// Retrieval info: PRIVATE: B_ACLR_SRC_MULT0 NUMERIC "3"
// Retrieval info: PRIVATE: B_CLK_SRC_MULT0 NUMERIC "0"
// Retrieval info: PRIVATE: CHAINOUT_OUTPUT_ACLR NUMERIC "3"
// Retrieval info: PRIVATE: CHAINOUT_OUTPUT_REG STRING "0"
// Retrieval info: PRIVATE: CHAINOUT_OUTPUT_REGISTER NUMERIC "0"
// Retrieval info: PRIVATE: CHAINOUT_OUTPUT_REGISTERED NUMERIC "0"
// Retrieval info: PRIVATE: CHAS_ZERO_CHAINOUT NUMERIC "0"
// Retrieval info: PRIVATE: EXTRA_MULTIPLIER_LATENCY NUMERIC "0"
// Retrieval info: PRIVATE: HAS_ACCUMULATOR NUMERIC "1"
// Retrieval info: PRIVATE: HAS_ACUMM_SLOAD NUMERIC "0"
// Retrieval info: PRIVATE: HAS_CHAININ_PORT NUMERIC "0"
// Retrieval info: PRIVATE: HAS_CHAINOUT_ADDER NUMERIC "0"
// Retrieval info: PRIVATE: HAS_LOOPBACK NUMERIC "0"
// Retrieval info: PRIVATE: HAS_MAC STRING "1"
// Retrieval info: PRIVATE: HAS_SAT_ROUND STRING "0"
// Retrieval info: PRIVATE: HAS_ZERO_LOOPBACK NUMERIC "0"
// Retrieval info: PRIVATE: IMPL_STYLE_DEDICATED NUMERIC "0"
// Retrieval info: PRIVATE: IMPL_STYLE_DEFAULT NUMERIC "1"
// Retrieval info: PRIVATE: IMPL_STYLE_LCELL NUMERIC "0"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix III"
// Retrieval info: PRIVATE: MULT_LATENCY NUMERIC "0"
// Retrieval info: PRIVATE: MULT_REGA0 NUMERIC "1"
// Retrieval info: PRIVATE: MULT_REGB0 NUMERIC "1"
// Retrieval info: PRIVATE: MULT_REGOUT0 NUMERIC "1"
// Retrieval info: PRIVATE: NUM_MULT STRING "2"
// Retrieval info: PRIVATE: OP1 STRING "Add"
// Retrieval info: PRIVATE: OP3 STRING "Add"
// Retrieval info: PRIVATE: OUTPUT_EXTRA_LAT NUMERIC "0"
// Retrieval info: PRIVATE: OUTPUT_REG_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: OUTPUT_REG_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: OVERFLOW NUMERIC "0"
// Retrieval info: PRIVATE: Q_ACLR_SRC_MULT0 NUMERIC "3"
// Retrieval info: PRIVATE: Q_CLK_SRC_MULT0 NUMERIC "0"
// Retrieval info: PRIVATE: REG_OUT NUMERIC "1"
// Retrieval info: PRIVATE: RNFORMAT STRING "44"
// Retrieval info: PRIVATE: ROTATE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ROTATE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ROTATE_OUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ROTATE_OUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ROTATE_OUT_REG STRING "1"
// Retrieval info: PRIVATE: ROTATE_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ROTATE_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ROTATE_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: ROTATE_REG STRING "1"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_MODE STRING "Disabled"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_OUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_OUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_OUT_REG STRING "0"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: ROUND3_CHAINOUT_REG STRING "1"
// Retrieval info: PRIVATE: ROUND3_FRAC_WIDTH NUMERIC "23"
// Retrieval info: PRIVATE: ROUND3_OUTPUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ROUND3_OUTPUT_CHAINOUT_TYPE STRING "Nearest Integer"
// Retrieval info: PRIVATE: ROUND3_OUTPUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ROUND3_OUTPUT_MODE STRING "Disabled"
// Retrieval info: PRIVATE: ROUND3_OUTPUT_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ROUND3_OUTPUT_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ROUND3_OUTPUT_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: ROUND3_OUTPUT_REG STRING "1"
// Retrieval info: PRIVATE: RQFORMAT STRING "Q1.30"
// Retrieval info: PRIVATE: RTS_WIDTH STRING "44"
// Retrieval info: PRIVATE: SAME_CONFIG NUMERIC "1"
// Retrieval info: PRIVATE: SAME_CONTROL_SRC_A0 NUMERIC "1"
// Retrieval info: PRIVATE: SAME_CONTROL_SRC_B0 NUMERIC "1"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_MODE STRING "Enabled"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_OUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_OUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: SAT3_CHAINOUT_REG STRING "1"
// Retrieval info: PRIVATE: SAT3_FRAC_WIDTH NUMERIC "1"
// Retrieval info: PRIVATE: SAT3_OUTPUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SAT3_OUTPUT_CHAINOUT_TYPE STRING "Symmetric"
// Retrieval info: PRIVATE: SAT3_OUTPUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SAT3_OUTPUT_MODE STRING "Enabled"
// Retrieval info: PRIVATE: SAT3_OUTPUT_OVERFLOW NUMERIC "0"
// Retrieval info: PRIVATE: SAT3_OUTPUT_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SAT3_OUTPUT_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SAT3_OUTPUT_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: SAT3_OUTPUT_REG STRING "1"
// Retrieval info: PRIVATE: SCANOUTA NUMERIC "0"
// Retrieval info: PRIVATE: SCANOUTB NUMERIC "0"
// Retrieval info: PRIVATE: SHIFTOUTA_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SHIFTOUTA_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SHIFTOUTA_REG STRING "0"
// Retrieval info: PRIVATE: SHIFT_RIGHT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SHIFT_RIGHT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SHIFT_RIGHT_OUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SHIFT_RIGHT_OUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SHIFT_RIGHT_OUT_REG STRING "1"
// Retrieval info: PRIVATE: SHIFT_RIGHT_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SHIFT_RIGHT_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SHIFT_RIGHT_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: SHIFT_RIGHT_REG STRING "1"
// Retrieval info: PRIVATE: SHIFT_ROTATE_MODE STRING "None"
// Retrieval info: PRIVATE: SIGNA STRING "SIGNED"
// Retrieval info: PRIVATE: SIGNA_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SIGNA_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SIGNA_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SIGNA_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SIGNA_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: SIGNA_REG STRING "1"
// Retrieval info: PRIVATE: SIGNB STRING "SIGNED"
// Retrieval info: PRIVATE: SIGNB_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SIGNB_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SIGNB_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SIGNB_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SIGNB_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: SIGNB_REG STRING "1"
// Retrieval info: PRIVATE: SRCA0 STRING "Multiplier input"
// Retrieval info: PRIVATE: SRCB0 STRING "Multiplier input"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: WIDTHA STRING "16"
// Retrieval info: PRIVATE: WIDTHB STRING "16"
// Retrieval info: PRIVATE: WIDTH_UPPER_DATA NUMERIC "1"
// Retrieval info: PRIVATE: ZERO_CHAINOUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ZERO_CHAINOUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ZERO_CHAINOUT_REG STRING "0"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_OUT_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_OUT_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_OUT_REG STRING "1"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: ZERO_LOOPBACK_REG STRING "1"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: ACCUMULATOR STRING "YES"
// Retrieval info: CONSTANT: ACCUM_DIRECTION STRING "ADD"
// Retrieval info: CONSTANT: ACCUM_SLOAD_ACLR STRING "ACLR3"
// Retrieval info: CONSTANT: ACCUM_SLOAD_PIPELINE_ACLR STRING "ACLR3"
// Retrieval info: CONSTANT: ACCUM_SLOAD_PIPELINE_REGISTER STRING "CLOCK0"
// Retrieval info: CONSTANT: ACCUM_SLOAD_REGISTER STRING "CLOCK0"
// Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_ACLR1 STRING "ACLR3"
// Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_PIPELINE_ACLR1 STRING "ACLR3"
// Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_PIPELINE_REGISTER1 STRING "CLOCK0"
// Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_REGISTER1 STRING "CLOCK0"
// Retrieval info: CONSTANT: CHAINOUT_ADDER STRING "NO"
// Retrieval info: CONSTANT: CHAINOUT_REGISTER STRING "UNREGISTERED"
// Retrieval info: CONSTANT: DEDICATED_MULTIPLIER_CIRCUITRY STRING "AUTO"
// Retrieval info: CONSTANT: INPUT_ACLR_A0 STRING "ACLR3"
// Retrieval info: CONSTANT: INPUT_ACLR_A1 STRING "ACLR3"
// Retrieval info: CONSTANT: INPUT_ACLR_B0 STRING "ACLR3"
// Retrieval info: CONSTANT: INPUT_ACLR_B1 STRING "ACLR3"
// Retrieval info: CONSTANT: INPUT_REGISTER_A0 STRING "CLOCK0"
// Retrieval info: CONSTANT: INPUT_REGISTER_A1 STRING "CLOCK0"
// Retrieval info: CONSTANT: INPUT_REGISTER_B0 STRING "CLOCK0"
// Retrieval info: CONSTANT: INPUT_REGISTER_B1 STRING "CLOCK0"
// Retrieval info: CONSTANT: INPUT_SOURCE_A0 STRING "DATAA"
// Retrieval info: CONSTANT: INPUT_SOURCE_A1 STRING "DATAA"
// Retrieval info: CONSTANT: INPUT_SOURCE_B0 STRING "DATAB"
// Retrieval info: CONSTANT: INPUT_SOURCE_B1 STRING "DATAB"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix III"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altmult_add"
// Retrieval info: CONSTANT: MULTIPLIER1_DIRECTION STRING "ADD"
// Retrieval info: CONSTANT: MULTIPLIER_ACLR0 STRING "ACLR3"
// Retrieval info: CONSTANT: MULTIPLIER_ACLR1 STRING "ACLR3"
// Retrieval info: CONSTANT: MULTIPLIER_REGISTER0 STRING "CLOCK0"
// Retrieval info: CONSTANT: MULTIPLIER_REGISTER1 STRING "CLOCK0"
// Retrieval info: CONSTANT: NUMBER_OF_MULTIPLIERS NUMERIC "2"
// Retrieval info: CONSTANT: OUTPUT_ACLR STRING "ACLR3"
// Retrieval info: CONSTANT: OUTPUT_REGISTER STRING "CLOCK0"
// Retrieval info: CONSTANT: PORT_ADDNSUB1 STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_SIGNA STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_SIGNB STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: REPRESENTATION_A STRING "SIGNED"
// Retrieval info: CONSTANT: REPRESENTATION_B STRING "SIGNED"
// Retrieval info: CONSTANT: SIGNED_ACLR_A STRING "ACLR3"
// Retrieval info: CONSTANT: SIGNED_ACLR_B STRING "ACLR3"
// Retrieval info: CONSTANT: SIGNED_PIPELINE_ACLR_A STRING "ACLR3"
// Retrieval info: CONSTANT: SIGNED_PIPELINE_ACLR_B STRING "ACLR3"
// Retrieval info: CONSTANT: SIGNED_PIPELINE_REGISTER_A STRING "CLOCK0"
// Retrieval info: CONSTANT: SIGNED_PIPELINE_REGISTER_B STRING "CLOCK0"
// Retrieval info: CONSTANT: SIGNED_REGISTER_A STRING "CLOCK0"
// Retrieval info: CONSTANT: SIGNED_REGISTER_B STRING "CLOCK0"
// Retrieval info: CONSTANT: WIDTH_A NUMERIC "16"
// Retrieval info: CONSTANT: WIDTH_B NUMERIC "16"
// Retrieval info: CONSTANT: WIDTH_CHAININ NUMERIC "1"
// Retrieval info: CONSTANT: WIDTH_RESULT NUMERIC "44"
// Retrieval info: CONSTANT: ZERO_CHAINOUT_OUTPUT_REGISTER STRING "UNREGISTERED"
// Retrieval info: CONSTANT: ZERO_LOOPBACK_ACLR STRING "ACLR3"
// Retrieval info: CONSTANT: ZERO_LOOPBACK_OUTPUT_ACLR STRING "ACLR3"
// Retrieval info: CONSTANT: ZERO_LOOPBACK_OUTPUT_REGISTER STRING "CLOCK0"
// Retrieval info: CONSTANT: ZERO_LOOPBACK_PIPELINE_ACLR STRING "ACLR3"
// Retrieval info: CONSTANT: ZERO_LOOPBACK_PIPELINE_REGISTER STRING "CLOCK0"
// Retrieval info: CONSTANT: ZERO_LOOPBACK_REGISTER STRING "CLOCK0"
// Retrieval info: USED_PORT: accum_sload 0 0 0 0 INPUT GND "accum_sload"
// Retrieval info: USED_PORT: aclr3 0 0 0 0 INPUT GND "aclr3"
// Retrieval info: USED_PORT: clock0 0 0 0 0 INPUT VCC "clock0"
// Retrieval info: USED_PORT: dataa_0 0 0 16 0 INPUT GND "dataa_0[15..0]"
// Retrieval info: USED_PORT: dataa_1 0 0 16 0 INPUT GND "dataa_1[15..0]"
// Retrieval info: USED_PORT: datab_0 0 0 16 0 INPUT GND "datab_0[15..0]"
// Retrieval info: USED_PORT: datab_1 0 0 16 0 INPUT GND "datab_1[15..0]"
// Retrieval info: USED_PORT: ena0 0 0 0 0 INPUT VCC "ena0"
// Retrieval info: USED_PORT: result 0 0 44 0 OUTPUT GND "result[43..0]"
// Retrieval info: CONNECT: @accum_sload 0 0 0 0 accum_sload 0 0 0 0
// Retrieval info: CONNECT: @aclr3 0 0 0 0 aclr3 0 0 0 0
// Retrieval info: CONNECT: @clock0 0 0 0 0 clock0 0 0 0 0
// Retrieval info: CONNECT: @dataa 0 0 16 0 dataa_0 0 0 16 0
// Retrieval info: CONNECT: @dataa 0 0 16 16 dataa_1 0 0 16 0
// Retrieval info: CONNECT: @datab 0 0 16 0 datab_0 0 0 16 0
// Retrieval info: CONNECT: @datab 0 0 16 16 datab_1 0 0 16 0
// Retrieval info: CONNECT: @ena0 0 0 0 0 ena0 0 0 0 0
// Retrieval info: CONNECT: result 0 0 44 0 @result 0 0 44 0
// Retrieval info: GEN_FILE: TYPE_NORMAL mult.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL mult.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mult.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mult.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mult_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mult_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf



