	
`define LAYER1_IN_FEATURE_ADDR_WIDTH 10
`define LAYER2_IN_FEATURE_ADDR_WIDTH 9
`define LAYER3_IN_FEATURE_ADDR_WIDTH 9
`define LAYER4_IN_FEATURE_ADDR_WIDTH 9

`define DATA_WIDTH 16
`define LAYER1_NUM_MULT 5
`define LAYER2_NUM_MULT 25

`define LAYER3_PO 25
`define LAYER4_PO 1