	
`define LAYER1_IN_FEATURE_ADDR_WIDTH 10
`define LAYER2_IN_FEATURE_ADDR_WIDTH 9
`define LAYER3_IN_FEATURE_ADDR_WIDTH 9


`define DATA_WIDTH 16
`define LAYER1_NUM_MULT 10
`define LAYER2_NUM_MULT 25
  

`define LAYER3_PO 4