`define LAYER1_IN_FEATURE_ADDR_WIDTH 10
`define LAYER2_IN_FEATURE_ADDR_WIDTH 9
`define LAYER3_IN_FEATURE_ADDR_WIDTH 9
`define LAYER4_IN_FEATURE_ADDR_WIDTH 9
`define LAYER5_IN_FEATURE_ADDR_WIDTH 9

`define DATA_WIDTH 16
`define LAYER1_NUM_MULT 20
`define LAYER2_NUM_MULT 20
`define LAYER3_NUM_MULT 2
`define LAYER3_NUM_MULT 20
`define IN_FEATURE_ADDR_WIDTH 10

`define INPUT_NUM_MEM  1  


`define LAYER4_PO 4