	
`define LAYER1_IN_FEATURE_ADDR_WIDTH 12
`define LAYER2_IN_FEATURE_ADDR_WIDTH 11
`define LAYER3_IN_FEATURE_ADDR_WIDTH 9
`define LAYER4_IN_FEATURE_ADDR_WIDTH 9

`define DATA_WIDTH 16
`define LAYER1_NUM_MULT 3
`define LAYER2_NUM_MULT 3

`define LAYER3_PO 2
`define LAYER4_PO 1